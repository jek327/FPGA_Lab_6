`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/22/2025 06:47:12 PM
// Design Name: 
// Module Name: D_FF_A
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module D_FF_A(input d, rstn, clk, output reg q);
    always @(posedge clk or negedge rstn)
    if (!rstn)
        q <= 0;
    else
        q <= d;
endmodule
